----------------------------------------------------------------------
-- @file    ENTITY_NAME.vhd
-- @brief   Entity implementation for ENTITY_NAME
-- @date    DATE_CREATED
-- @version v1.0.0
-- @author  AUTHORS
----------------------------------------------------------------------

------ LIBRARY & USE STATEMENTS ------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--------- ENTITY DECLARATION ---------
entity ENTITY_NAME is
    generic (
        --! Define generic properties here
    );
    port (
        --! Define inputs/outputs here
    );
end ENTITY_NAME;

------ Architecture Declaration ------
architecture rtl of ENTITY_NAME is
    ------------ COMPONENTS --------------
    --! Add component definitions here

    -------------- SIGNALS ---------------
    --! Add internal signals here

    ------------- CONSTANTS --------------
    --! Add constants here
begin
    --! Implement your entity here
end rtl;